module top (
    input wire clk, // 50mhz clock
    input wire [3:0] btn,
    input wire [9:0] sw,
    input wire uart_rx,
    output wire uart_tx,
    output wire [9:0] led
);



    
endmodule
