module top (
    input wire clk,
    input wire reset,
    input wire rx,
    output wire tx,
    output wire [3:0]led,
    inout [13:0]ck_io
);


always @(posedge clk) begin

end

endmodule
